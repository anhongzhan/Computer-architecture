`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:44:57 10/19/2018
// Design Name:   alu
// Module Name:   F:/ise project/alu/alu_test.v
// Project Name:  alu
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: alu
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module alu_test;

	// Inputs
	reg [31:0] A;
	reg [31:0] B;
	reg [4:0] Card;
	reg Cin;

	// Outputs
	wire [31:0] F;
	wire Cout;
	wire Zero;

	// Instantiate the Unit Under Test (UUT)
	alu uut (
		.A(A), 
		.B(B), 
		.Card(Card), 
		.Cin(Cin), 
		.F(F), 
		.Cout(Cout), 
		.Zero(Zero)
	);

	initial begin
		// Initialize Inputs
		A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b00001;
		Cin = 0;

		// Wait 10 ns for global reset to finish
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b00010;
		Cin = 0;  
		// Add stimulus here
		#10;
		A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b00011;
		Cin = 0; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b00100;
		Cin = 0; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b00101;
		Cin = 0; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b00110;
		Cin = 0; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b00111;
		Cin = 0; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01000;
		Cin = 0; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01001;
		Cin = 1; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01010;
		Cin = 1; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01011;
		Cin = 1; 
		
		#10;
		A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01100;
		Cin = 1;
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01101;
		Cin = 1; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01110;
		Cin = 1; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b01111;
		Cin = 1; 
		
		#10;
      A = 32'b10101010101010101010101010101010;
		B = 32'b11001100110011001100110011001100;
		Card = 5'b10000;
		Cin = 1; 
		
		#10;
	end
      
endmodule

